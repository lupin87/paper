 //date:16/11/2011
`timescale 1ns/1ps
//`include "./test_core.v"
// `include "./test_core_new.v"
//`include "./test_core_new.v"
module test_core_tb;

//khai bao bien ngo vao
reg clk;
reg start;
reg reset;
//reg [7:0]fram_datain;

//khai bao bien ngo ra
wire result_ack;//bao ket thuc nhan dang
wire [5:0]result;//chi so tu
wire overflow;//bao ket qua nhan dang khong dang tin cay

//goi module test
test_core test_core(result_ack,result,overflow,start,clk,reset);
`include "./dump.v"

//  initial
//      begin
//	 #30000ns $finish;
//       end
initial begin
     $vcdpluson(1,test_core_tb);
     $vcdpluson(0,test_core_tb.test_core);
end // initial begin

integer f;
always @ (result_ack)
      begin
       if (result_ack == 1'b1) begin
        f = $fopen("output.txt");
        $fmonitor(f, "time=%5d, result=%d\n", $time,result[5:0] );
        $display("time=%5d, result=%d\n", $time,result[5:0] );
        #500;
        $fclose(f);
        $finish;
       end
      end // initial begin
////gan gia tri ngo vao
initial
begin
 clk=1'b0;
 reset=1'b0;
 start=1'b0;
 //fram_datain=0;//from Speech RAM
 #20
 reset=1'b1;
 start=1'b0;
 $display ("data_in = %h", test_core.fecore.ram_datain);
 /*
 #120
 fram_datain=2;
 #20//bat dau subframe 1
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20//ket thuc subframe 1
 fram_datain=10;
 
 #20//8 bit thap cua mau thu nhat subframe 2, t=3270
 fram_datain=2;
 

 #53600//subframe 2 (tiep 8 bit cao cua mau thu nhat va doc tiep cac mau con lai), t=56870
 fram_datain=4;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=-5;
 #20
 fram_datain=-10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=45;
 #20
 fram_datain=76;
 #20
 fram_datain=-23;
 #20
 fram_datain=10;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=85;
 #20
 fram_datain=24;
 #20
 fram_datain=5;
 #20
 fram_datain=2;
 #20
 fram_datain=80;
 #20
 fram_datain=27;
 #20
 fram_datain=30;
 #20
 fram_datain=40;
 #20
 fram_datain=15;
 #20
 fram_datain=36;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=4;
 #20
 fram_datain=21;
 #20
 fram_datain=16;
 #20
 fram_datain=18;
 #20
 fram_datain=32;
 #20
 fram_datain=9;
 #20
 fram_datain=35;
 #20
 fram_datain=100;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=105;
 #20
 fram_datain=115;
 #20
 fram_datain=120;
 #20
 fram_datain=125;
 #20
 fram_datain=130;
 #20
 fram_datain=135;
 #20
 fram_datain=140;
 #20
 fram_datain=145;
 #20
 fram_datain=150;
 #20
 fram_datain=155;
 #20
 fram_datain=-5;
 #20
 fram_datain=-10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=45;
 #20
 fram_datain=76;
 #20
 fram_datain=-23;
 #20
 fram_datain=10;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=85;
 #20
 fram_datain=24;
 
 #20//bat dau subframe 3
 fram_datain=5;
 
 #53600//t=113650
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=5;
 #20
 fram_datain=10;
 #20
 fram_datain=15;
 #20
 fram_datain=20;
 #20
 fram_datain=25;
 #20
 fram_datain=30;
 #20
 fram_datain=35;
 #20
 fram_datain=40;
 #20
 fram_datain=45;
 #20
 fram_datain=50;
 #20
 fram_datain=55;
 #20
 fram_datain=60;
 #20
 fram_datain=65;
 #20
 fram_datain=70;
 #20
 fram_datain=75;
 #20
 fram_datain=80;
 #20
 fram_datain=85;
 #20
 fram_datain=90;
 #20
 fram_datain=95;
 #20
 fram_datain=100;
 #20
 fram_datain=0;
 #20//ket thuc subframe 3
 fram_datain=0;
 
 #20//bat dau subframe 4
 fram_datain=0;
 
 #53600//t=170430
 fram_datain=0;
 #20
 fram_datain=0;
 */
 end
 always
 #10
 clk=~clk;
 endmodule


